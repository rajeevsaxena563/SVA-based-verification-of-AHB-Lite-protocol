`include "definesPkg.sv"
`include "AHB_interface.sv"
`include "ahb_generator.sv"
`include "ahb_driver.sv"
`include "ahb_environment.sv"
`include "ahbSlave.sv"
`include "AHBSlave_top.sv"
`include "ahb_test.sv"
`include "ahb_top.sv"
`include "assertions.sv"
